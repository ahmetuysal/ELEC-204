library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

entity SEVSEG_CLOCK_GENERATOR is
    Port ( MCLK : in  STD_LOGIC;
           SEVSEG_CLOCK : out  STD_LOGIC);
end SEVSEG_CLOCK_GENERATOR;

architecture Behavioral of SEVSEG_CLOCK_GENERATOR is

SIGNAL COUNTER: STD_LOGIC_VECTOR(17 DOWNTO 0) := "000000000000000000";

begin

PROCESS(MCLK)

BEGIN

	IF(MCLK'EVENT AND MCLK = '1') THEN
		IF COUNTER < "101101110001101100" THEN
			COUNTER <= COUNTER + 1;
		ELSE
			COUNTER <= "000000000000000000";
		END IF;
	END IF;
END PROCESS;

SEVSEG_CLOCK <= '1' WHEN COUNTER < "010110111000110110"
ELSE '0';


end Behavioral;

