----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    14:46:24 11/17/2017 
-- Design Name: 
-- Module Name:    SEVSEG_DRIVER - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity SEVSEG_DRIVER is
    Port ( C1 : in  STD_LOGIC_VECTOR (10 downto 0);
           C2 : in  STD_LOGIC_VECTOR (10 downto 0);
           C3 : in  STD_LOGIC_VECTOR (10 downto 0);
           C4 : in  STD_LOGIC_VECTOR (10 downto 0);
           CLK : in  STD_LOGIC;
			  SELECTING_DISPLAY_INPUT : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
			  ISSELECTING : IN STD_LOGIC;
			  SELECT_COUNTER : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
           SEVSEG_DATA_BCD : out  STD_LOGIC_VECTOR (3 downto 0);
           SEVSEG_DRIVER : out  STD_LOGIC_VECTOR (7 downto 0));
end SEVSEG_DRIVER;

architecture Behavioral of SEVSEG_DRIVER is

SIGNAL COUNTER : STD_LOGIC_VECTOR(2 DOWNTO 0) := "000";
SIGNAL SELECTING_BCD_1 : STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL SELECTING_BCD_2 : STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL DISPLAYING_BCD : STD_LOGIC_VECTOR(15 DOWNTO 0);
-- PROCEDURE DENEME --
-- DOUBLE DABBLE ALGORITHM --
PROCEDURE F_5BIT_BINARY_2_8BIT_BCD (
	SIGNAL FIVEBIT_BINARY_IN : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
	SIGNAL RESULT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	)IS
		
		VARIABLE TEMP : STD_LOGIC_VECTOR(4 DOWNTO 0);
		VARIABLE BCD : UNSIGNED(7 DOWNTO 0);
		
		BEGIN
		--Zero the bcd var
		BCD := (OTHERS => '0');
		--Read input to temp var
		TEMP(4 DOWNTO 0) := FIVEBIT_BINARY_IN;
		
		--Cycle 5 times (number of input bits)
		
		FOR I IN 0 TO 4 LOOP
		
			IF(BCD(3 DOWNTO 0) >  4) THEN
				BCD(3 DOWNTO 0) := BCD(3 DOWNTO 0) +3;
			END IF;
			--shift bcd left 1 bit, concatanate with msb of temp
			BCD := BCD(6 DOWNTO 0) & TEMP(4);
			--Shift temp left 1 bit
			TEMP := TEMP(3 DOWNTO 0) & '0';
		END LOOP;
			
		RESULT <= STD_LOGIC_VECTOR(BCD);
			
END PROCEDURE F_5BIT_BINARY_2_8BIT_BCD;

PROCEDURE F_11BIT_BINARY_2_16BIT_BCD (
	SIGNAL ELEVENBIT_BINARY_IN : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
	SIGNAL RESULT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	)IS
		
		VARIABLE TEMP : STD_LOGIC_VECTOR(10 DOWNTO 0);
		VARIABLE BCD : UNSIGNED(15 DOWNTO 0);
		
		BEGIN
		--Zero the bcd var
		BCD := (OTHERS => '0');
		--Read input to temp var
		TEMP(10 DOWNTO 0) := ELEVENBIT_BINARY_IN;
		
		--Cycle 11 times (number of input bits)
		
		FOR I IN 0 TO 10 LOOP
		
			IF(BCD(3 DOWNTO 0) >  4) THEN
				BCD(3 DOWNTO 0) := BCD(3 DOWNTO 0) +3;
			END IF;
			
			IF(BCD(7 DOWNTO 4) > 4) THEN
				BCD(7 DOWNTO 4) := BCD(7 DOWNTO 4)+3;
			END IF;
			
			IF(BCD(11 DOWNTO 8) > 4) THEN
				BCD(11 DOWNTO 8) := BCD(11 DOWNTO 8)+3;
			END IF;
			--shift bcd left 1 bit, concatanate with msb of temp
			BCD := BCD(14 DOWNTO 0) & TEMP(10);
			--Shift temp left 1 bit
			TEMP := TEMP(9 DOWNTO 0) & '0';
		END LOOP;
			
		RESULT <= STD_LOGIC_VECTOR(BCD);
			
END PROCEDURE F_11BIT_BINARY_2_16BIT_BCD;

-- PROCEDURE DENEME --
begin

	PROCESS_CLK : PROCESS(CLK)
	BEGIN 
		IF (CLK'EVENT AND CLK = '1') THEN
			COUNTER <= COUNTER +1 ;
		END IF;
	END PROCESS;
	
	-- SELECTING SEVSEG CELL TO UPDATE 
	WITH COUNTER SELECT SEVSEG_DRIVER <=
	"01111111" WHEN "000",
	"10111111" WHEN "001",
	"11011111" WHEN "010",
	"11101111" WHEN "011",
	"11110111" WHEN "100",
	"11111011" WHEN "101",
	"11111101" WHEN "110",
	"11111110" WHEN "111",
	"00001111" WHEN OTHERS;

	-- SELECTING SEVSEG DATA TO DISPLAY 
	PROCESS(ISSELECTING,SELECT_COUNTER,SELECTING_DISPLAY_INPUT,COUNTER,C1,C2,C3,C4)
		BEGIN
		IF (ISSELECTING = '1') THEN --WE ARE ON SELECTION PHASE
			IF(SELECT_COUNTER = "00") THEN -- WE ARE SELECTING A1 AND A2
			F_5BIT_BINARY_2_8BIT_BCD(SELECTING_DISPLAY_INPUT(9 DOWNTO 5),SELECTING_BCD_1);
			F_5BIT_BINARY_2_8BIT_BCD(SELECTING_DISPLAY_INPUT(4 DOWNTO 0),SELECTING_BCD_2);
			CASE(COUNTER) IS 
			WHEN "000" => 
				SEVSEG_DATA_BCD <= "1010"; --A
			WHEN "001" => 
				SEVSEG_DATA_BCD <= "0001"; --1
			WHEN "010" => 
				SEVSEG_DATA_BCD <= SELECTING_BCD_1(7 DOWNTO 4);
			WHEN "011" => 
				SEVSEG_DATA_BCD <= SELECTING_BCD_1(3 DOWNTO 0);
			WHEN "100" => 
				SEVSEG_DATA_BCD <= "1010"; --A
			WHEN "101" => 
				SEVSEG_DATA_BCD <= "0010"; --2
			WHEN "110" => 
				SEVSEG_DATA_BCD <= SELECTING_BCD_2(7 DOWNTO 4);
			WHEN "111" => 
				SEVSEG_DATA_BCD <= SELECTING_BCD_2(3 DOWNTO 0);
			WHEN OTHERS => 
				NULL;
			END CASE;
			ELSIF(SELECT_COUNTER = "01") THEN -- SELECTING A3,A4
			F_5BIT_BINARY_2_8BIT_BCD(SELECTING_DISPLAY_INPUT(9 DOWNTO 5),SELECTING_BCD_1);
			F_5BIT_BINARY_2_8BIT_BCD(SELECTING_DISPLAY_INPUT(4 DOWNTO 0),SELECTING_BCD_2);
			CASE(COUNTER) IS 
			WHEN "000" => 
				SEVSEG_DATA_BCD <= "1010"; --A
			WHEN "001" => 
				SEVSEG_DATA_BCD <= "0011"; --3
			WHEN "010" => 
				SEVSEG_DATA_BCD <= SELECTING_BCD_1(7 DOWNTO 4);
			WHEN "011" => 
				SEVSEG_DATA_BCD <= SELECTING_BCD_1(3 DOWNTO 0);
			WHEN "100" => 
				SEVSEG_DATA_BCD <= "1010"; --A
			WHEN "101" => 
				SEVSEG_DATA_BCD <= "0100"; --4
			WHEN "110" => 
				SEVSEG_DATA_BCD <= SELECTING_BCD_2(7 DOWNTO 4);
			WHEN "111" => 
				SEVSEG_DATA_BCD <= SELECTING_BCD_2(3 DOWNTO 0);
			WHEN OTHERS => 
				NULL;
			END CASE;
			ELSIF(SELECT_COUNTER = "10") THEN -- SELECTING B1,B2
				F_5BIT_BINARY_2_8BIT_BCD(SELECTING_DISPLAY_INPUT(9 DOWNTO 5),SELECTING_BCD_1);
				F_5BIT_BINARY_2_8BIT_BCD(SELECTING_DISPLAY_INPUT(4 DOWNTO 0),SELECTING_BCD_2);
				CASE(COUNTER) IS 
				WHEN "000" => 
					SEVSEG_DATA_BCD <= "1011"; --B
				WHEN "001" => 
					SEVSEG_DATA_BCD <= "0001"; --1
				WHEN "010" => 
					SEVSEG_DATA_BCD <= SELECTING_BCD_1(7 DOWNTO 4);
				WHEN "011" => 
					SEVSEG_DATA_BCD <= SELECTING_BCD_1(3 DOWNTO 0);
				WHEN "100" => 
					SEVSEG_DATA_BCD <= "1011"; --B
				WHEN "101" => 
					SEVSEG_DATA_BCD <= "0010"; --2
				WHEN "110" => 
					SEVSEG_DATA_BCD <= SELECTING_BCD_2(7 DOWNTO 4);
				WHEN "111" => 
					SEVSEG_DATA_BCD <= SELECTING_BCD_2(3 DOWNTO 0);
				WHEN OTHERS => 
					NULL;
				END CASE;
			ELSIF(SELECT_COUNTER = "11") THEN -- SELECTING B3,B4
				F_5BIT_BINARY_2_8BIT_BCD(SELECTING_DISPLAY_INPUT(9 DOWNTO 5),SELECTING_BCD_1);
				F_5BIT_BINARY_2_8BIT_BCD(SELECTING_DISPLAY_INPUT(4 DOWNTO 0),SELECTING_BCD_2);
				CASE(COUNTER) IS 
				WHEN "000" => 
					SEVSEG_DATA_BCD <= "1011"; --B
				WHEN "001" => 
					SEVSEG_DATA_BCD <= "0011"; --3
				WHEN "010" => 
					SEVSEG_DATA_BCD <= SELECTING_BCD_1(7 DOWNTO 4);
				WHEN "011" => 
					SEVSEG_DATA_BCD <= SELECTING_BCD_1(3 DOWNTO 0);
				WHEN "100" => 
					SEVSEG_DATA_BCD <= "1011"; --B
				WHEN "101" => 
					SEVSEG_DATA_BCD <= "0100"; --4
				WHEN "110" => 
					SEVSEG_DATA_BCD <= SELECTING_BCD_2(7 DOWNTO 4);
				WHEN "111" => 
					SEVSEG_DATA_BCD <= SELECTING_BCD_2(3 DOWNTO 0);
				WHEN OTHERS => 
					NULL;
				END CASE;
			END IF;
		ELSE -- DISPLAYING THE RESULTS (2 RIGHTMOST SWITCHS ARE USED AS SELECTION INPUT) 
			IF(SELECTING_DISPLAY_INPUT(1 DOWNTO 0) = "00") THEN --DISPLAYING C1
				F_11BIT_BINARY_2_16BIT_BCD(C1,DISPLAYING_BCD);
				CASE(COUNTER) IS 
				WHEN "000" => 
					SEVSEG_DATA_BCD <= "1100"; --C
				WHEN "001" => 
					SEVSEG_DATA_BCD <= "0001"; --1
				WHEN "010" => 
					SEVSEG_DATA_BCD <= "1111"; --EMPTY
				WHEN "011" => 
					SEVSEG_DATA_BCD <= "1111"; --EMPTY
				WHEN "100" => 
					SEVSEG_DATA_BCD <= DISPLAYING_BCD(15 DOWNTO 12);
				WHEN "101" => 
					SEVSEG_DATA_BCD <= DISPLAYING_BCD(11 DOWNTO 8);
				WHEN "110" => 
					SEVSEG_DATA_BCD <= DISPLAYING_BCD(7 DOWNTO 4);
				WHEN "111" => 
					SEVSEG_DATA_BCD <= DISPLAYING_BCD(3 DOWNTO 0);
				WHEN OTHERS => 
					NULL;
				END CASE;
			ELSIF(SELECTING_DISPLAY_INPUT(1 DOWNTO 0) = "01") THEN -- DISPLAYING C2
				F_11BIT_BINARY_2_16BIT_BCD(C2,DISPLAYING_BCD);
				CASE(COUNTER) IS 
				WHEN "000" => 
					SEVSEG_DATA_BCD <= "1100"; --C
				WHEN "001" => 
					SEVSEG_DATA_BCD <= "0010"; --2
				WHEN "010" => 
					SEVSEG_DATA_BCD <= "1111"; --EMPTY
				WHEN "011" => 
					SEVSEG_DATA_BCD <= "1111"; --EMPTY
				WHEN "100" => 
					SEVSEG_DATA_BCD <= DISPLAYING_BCD(15 DOWNTO 12);
				WHEN "101" => 
					SEVSEG_DATA_BCD <= DISPLAYING_BCD(11 DOWNTO 8);
				WHEN "110" => 
					SEVSEG_DATA_BCD <= DISPLAYING_BCD(7 DOWNTO 4);
				WHEN "111" => 
					SEVSEG_DATA_BCD <= DISPLAYING_BCD(3 DOWNTO 0);
				WHEN OTHERS => 
					NULL;
				END CASE;
			ELSIF(SELECTING_DISPLAY_INPUT(1 DOWNTO 0) = "10") THEN -- DISPLAYING C3
				F_11BIT_BINARY_2_16BIT_BCD(C3,DISPLAYING_BCD);
				CASE(COUNTER) IS 
				WHEN "000" => 
					SEVSEG_DATA_BCD <= "1100"; --C
				WHEN "001" => 
					SEVSEG_DATA_BCD <= "0011"; --3
				WHEN "010" => 
					SEVSEG_DATA_BCD <= "1111"; --EMPTY
				WHEN "011" => 
					SEVSEG_DATA_BCD <= "1111"; --EMPTY
				WHEN "100" => 
					SEVSEG_DATA_BCD <= DISPLAYING_BCD(15 DOWNTO 12);
				WHEN "101" => 
					SEVSEG_DATA_BCD <= DISPLAYING_BCD(11 DOWNTO 8);
				WHEN "110" => 
					SEVSEG_DATA_BCD <= DISPLAYING_BCD(7 DOWNTO 4);
				WHEN "111" => 
					SEVSEG_DATA_BCD <= DISPLAYING_BCD(3 DOWNTO 0);
				WHEN OTHERS => 
					NULL;
				END CASE;
			ELSIF(SELECTING_DISPLAY_INPUT(1 DOWNTO 0) = "11") THEN -- DISPLAYING C4
				F_11BIT_BINARY_2_16BIT_BCD(C4,DISPLAYING_BCD);
				CASE(COUNTER) IS 
				WHEN "000" => 
					SEVSEG_DATA_BCD <= "1100"; --C
				WHEN "001" => 
					SEVSEG_DATA_BCD <= "0100"; --4
				WHEN "010" => 
					SEVSEG_DATA_BCD <= "1111"; --EMPTY
				WHEN "011" => 
					SEVSEG_DATA_BCD <= "1111"; --EMPTY
				WHEN "100" => 
					SEVSEG_DATA_BCD <= DISPLAYING_BCD(15 DOWNTO 12);
				WHEN "101" => 
					SEVSEG_DATA_BCD <= DISPLAYING_BCD(11 DOWNTO 8);
				WHEN "110" => 
					SEVSEG_DATA_BCD <= DISPLAYING_BCD(7 DOWNTO 4);
				WHEN "111" => 
					SEVSEG_DATA_BCD <= DISPLAYING_BCD(3 DOWNTO 0);
				WHEN OTHERS => 
					NULL;
				END CASE;
			END IF;
		END IF;
	END PROCESS;
end Behavioral;

